module not1bit (a,out);
    input a;
    output out;
    not(out,a);
endmodule