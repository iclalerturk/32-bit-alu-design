`include "alu.v"
module alu_tb;
    reg [31:0]a, b;
    reg [2:0]alu;
    wire [31:0]result;
    wire cout;
    

    alu add1(a,b,alu,result,cout);

    initial begin
        $dumpfile("alu.vcd");
        $dumpvars(0, alu_tb);
        a = 32'b00000000000000000000000011110000;
        b = 32'b00000000000000000000000000000001;
        alu = 3'b101;
        #1;
        a = 32'b10000000000000000000000011110000;
        b = 32'b00000000000000000000000000000001;
        alu = 3'b101;
        #1;
        a = 32'b00000000000000000000000011110000;
        b = 32'b00000000000000000000000000000001;
        alu = 3'b011;
        #1;
        a = 32'b00000000000000000000000011110000;
        b = 32'b00000000000000000000000000000001;
        alu = 3'b010;
        #1;
        a = 32'b00000000000000000000000011110000;
        b = 32'b00000000000000000000000000000001;
        alu = 3'b001;
        #1;
        a = 32'b00000000000000000000000011110000;
        b = 32'b00000000000000000000000000000001;
        alu = 3'b000;
        #1;
        //111:pass, 110:pass, 101:slt, 100:pass, 011:xor, 010:and, 001:sub, 000:sum
        //111:a, 110:b, 101:c, 100:d, 011:e, 010:f, 001:g, 000:h
    end
endmodule
//iverilog -o alu_tb.vvp alu_tb.v
//vvp alu_tb.vvp